module tb_full_adder;
reg a,b,cin;
wire sum,carry;

full_adder dut(a,b,cin,sum,carry);

initial begin
    $dumpfile("full_adder.vcd");
    $dumpvars(0, tb_full_adder);

    a=0;b=0;cin=0; #10;
    a=0;b=1;cin=0; #10;
    a=1;b=0;cin=1; #10;
    a=1;b=1;cin=1; #10;

    $finish;
end
endmodule
